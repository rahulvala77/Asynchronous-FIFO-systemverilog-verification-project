//-----------------------------------------------------------------------------------------------------------------------
//BLOCK - fifo_mem
//Description - It is queue array which can be used anywhere in ENV
//-----------------------------------------------------------------------------------------------------------------------

class fifo_mem;

  bit [7:0] queue[$];  //variable declaration => used in predicto,scoreboard

endclass
